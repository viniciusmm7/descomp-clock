tmp(0)	:= "0000000000000";	-- 	;COMENTARIO TESTE 1
tmp(1)	:= "0000000000000";	-- NOP 	;COMENTARIO TESTE 2
tmp(2)	:= "0001000000000";	-- LDA $0
tmp(3)	:= "0101100100000";	-- STA @288
tmp(4)	:= "0010000000001";	-- ADD $1
tmp(5)	:= "1100000000000";	-- AND 	;COMENTARIO TESTE 3
tmp(6)	:= "0110000000111";	-- JMP .TEST
tmp(7)	:= "0110000001000";	-- JMP .TEST2
tmp(8)	:= "1001000001010";	-- JSR .SUBROTINA_TESTE
tmp(9)	:= "0110000000111";	-- JMP .TEST
tmp(10)	:= "1000000000000";	-- RET 	;COMENTARIO TESTE 4
