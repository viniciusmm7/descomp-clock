tmp(0)	:= "0001000000000";	-- LDA $0
tmp(1)	:= "0101100100000";	-- STA @288
tmp(2)	:= "0010000000001";	-- ADD $1
tmp(3)	:= "0110000000100";	-- JMP .TEST
tmp(4)	:= "0110000000101";	-- JMP .TEST2
tmp(5)	:= "0110000000000";	-- JMP .LOOP
