tmp(0)	:= "0000000000000";	-- 	; SETUP
tmp(1)	:= "0101111111111";	-- STA @511    	; reseta a leitura do key 0
tmp(2)	:= "0101111111110";	-- STA @510    	; reseta a leitura do key 1
tmp(3)	:= "0101111111101";	-- STA @509    	; reseta a leitura do key reset
tmp(4)	:= "0100000000000";	-- LDI $0      	; carrega o valor inicial das casas
tmp(5)	:= "0101000111001";	-- STA @57     	; intervalo numérico de configuração
tmp(6)	:= "0101000000000";	-- STA @0      	; armazena 0 na unidade
tmp(7)	:= "0101000000001";	-- STA @1      	; armazena 0 na dezena
tmp(8)	:= "0101000000010";	-- STA @2      	; armazena 0 na centena
tmp(9)	:= "0101000000011";	-- STA @3      	; armazena 0 no milhar
tmp(10)	:= "0101000000100";	-- STA @4      	; armazena 0 na dezena de milhar
tmp(11)	:= "0101000000101";	-- STA @5      	; armazena 0 na centena de milhar
tmp(12)	:= "0101000001000";	-- STA @8      	; armazena um 0 de referência
tmp(13)	:= "0100000000001";	-- LDI $1      	; carrega o valor de incremento
tmp(14)	:= "0101000000110";	-- STA @6      	; armazena o valor de incremento
tmp(15)	:= "0101000001001";	-- STA @9			; armazena 1 no 9 para referência do intervalo numérico de configuração
tmp(16)	:= "0100000001010";	-- LDI $10     	; carrega o valor máximo por casa possível
tmp(17)	:= "0101000000111";	-- STA @7      	; armazena o valor máximo por casa possível
tmp(18)	:= "0100000001001";	-- LDI $9      	; carrega o número 9 para definir o limite de contagem inicial
tmp(19)	:= "0101000111010";	-- STA @58     	; armazena na casa das unidades do limite
tmp(20)	:= "0101000111011";	-- STA @59     	; armazena na casa das dezenas do limite
tmp(21)	:= "0101000111100";	-- STA @60     	; armazena na casa das centenas do limite
tmp(22)	:= "0101000111101";	-- STA @61     	; armazena na casa dos milhares do limite
tmp(23)	:= "0101000111110";	-- STA @62     	; armazena na casa das dezenas de milhar do limite
tmp(24)	:= "0101000111111";	-- STA @63     	; armazena na casa das centenas de milhar do limite
tmp(25)	:= "0100000000010";	-- LDI $2			; carrega 2 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(26)	:= "0101000001010";	-- STA @10			; armazena a referência de estado 2 no endereço 10
tmp(27)	:= "0100000000011";	-- LDI $3			; carrega 3 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(28)	:= "0101000001011";	-- STA @11			; armazena a referência de estado 3 no endereço 11
tmp(29)	:= "0100000000100";	-- LDI $4			; carrega 4 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(30)	:= "0101000001100";	-- STA @12			; armazena a referência de estado 4 no endereço 12
tmp(31)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(32)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(33)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(34)	:= "0111000100101";	-- JEQ .PULA_RESET
tmp(35)	:= "0101111111101";	-- STA @509
tmp(36)	:= "1001001001111";	-- JSR .RESET
tmp(37)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(38)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(39)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(40)	:= "0111000101011";	-- JEQ .PULA_CONFIG
tmp(41)	:= "0101111111110";	-- STA @510
tmp(42)	:= "0110000110111";	-- JMP .INICIO_LOOP_CONFIGURACAO_LIMITE
tmp(43)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(44)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(45)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(46)	:= "0111000110100";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(47)	:= "0101111111111";	-- STA @511
tmp(48)	:= "1001100111101";	-- JSR .ATINGIU_LIMITE			; verifica se a contagem atingiu o limite
tmp(49)	:= "1000000000110";	-- CEQ @6						; se atingiu o limite, pula o incrementa contagem
tmp(50)	:= "0111000110100";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(51)	:= "1001001010111";	-- JSR .INCREMENTA_CONTAGEM
tmp(52)	:= "1001011101111";	-- JSR .APAGA_LEDS         	; apaga os LEDs
tmp(53)	:= "1001010001000";	-- JSR .MOSTRA_CONTAGEM    	; escreve os números da contagem nos displays
tmp(54)	:= "0110000011111";	-- JMP .LOOP_PRINCIPAL
tmp(55)	:= "0100000000011";	-- LDI $3			; acende os leds da primeira posição
tmp(56)	:= "0101100000000";	-- STA @256
tmp(57)	:= "1001001001111";	-- JSR .RESET		; reseta a contagem
tmp(58)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(59)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(60)	:= "1000000000110";	-- CEQ @6      	; verifica se é 1
tmp(61)	:= "0111001001100";	-- JEQ .SAIR_LOOP_CONFIGURACAO_LIMITE
tmp(62)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(63)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(64)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(65)	:= "0111001000100";	-- JEQ .PULA_MUDANCA_ESTADO
tmp(66)	:= "0101111111110";	-- STA @510
tmp(67)	:= "0110001001100";	-- JMP .SAIR_LOOP_CONFIGURACAO_LIMITE
tmp(68)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(69)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(70)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(71)	:= "0111001001010";	-- JEQ .PULA_MUDANCA_INTERVALO
tmp(72)	:= "0101111111111";	-- STA @511
tmp(73)	:= "1001011110100";	-- JSR .MUDA_INTERVALO
tmp(74)	:= "1001010010101";	-- JSR .MOSTRA_LIMITE
tmp(75)	:= "0110000111010";	-- JMP .LOOP_CONFIGURACAO_LIMITE
tmp(76)	:= "0100000000000";	-- LDI $0    		; carrega 0
tmp(77)	:= "0101000111001";	-- STA @57     	; armazena 0 no intervalo de mudança atual
tmp(78)	:= "0110000011111";	-- JMP .LOOP_PRINCIPAL
tmp(79)	:= "0100000000000";	-- LDI $0
tmp(80)	:= "0101000000000";	-- STA @0
tmp(81)	:= "0101000000001";	-- STA @1
tmp(82)	:= "0101000000010";	-- STA @2
tmp(83)	:= "0101000000011";	-- STA @3
tmp(84)	:= "0101000000100";	-- STA @4
tmp(85)	:= "0101000000101";	-- STA @5
tmp(86)	:= "1010000000000";	-- RET
tmp(87)	:= "0001000000000";	-- LDA @0                  	; carrega o valor da unidade
tmp(88)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da unidade
tmp(89)	:= "1000000000111";	-- CEQ @7                  	; compara o valor da casa com 10
tmp(90)	:= "0111001011101";	-- JEQ .INCREMENTA_DEZENA  	; incrementa a casa da dezena caso necessário
tmp(91)	:= "0101000000000";	-- STA @0                  	; armazena o valor da unidade
tmp(92)	:= "1010000000000";	-- RET
tmp(93)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(94)	:= "0101000000000";	-- STA @0                  	; armazena 0 na unidade
tmp(95)	:= "0001000000001";	-- LDA @1                  	; carrega o valor atual da dezena
tmp(96)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena
tmp(97)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(98)	:= "0111001100101";	-- JEQ .INCREMENTA_CENTENA 	; se for, incrementa a centena
tmp(99)	:= "0101000000001";	-- STA @1                  	; armazena o novo valor da dezena
tmp(100)	:= "0110001011100";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(101)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(102)	:= "0101000000001";	-- STA @1                  	; armazena 0 na dezena
tmp(103)	:= "0001000000010";	-- LDA @2                  	; carrega o valor atual da centena
tmp(104)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena
tmp(105)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(106)	:= "0111001101101";	-- JEQ .INCREMENTA_MILHAR  	; se for, incrementa o milhar
tmp(107)	:= "0101000000010";	-- STA @2                  	; armazena o novo valor da centena
tmp(108)	:= "0110001011100";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(109)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(110)	:= "0101000000010";	-- STA @2                  	; armazena 0 na centena
tmp(111)	:= "0001000000011";	-- LDA @3                  	; carrega o valor atual do milhar
tmp(112)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor do milhar
tmp(113)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(114)	:= "0111001110101";	-- JEQ .INCREMENTA_DMILHAR 	; se for, incrementa a dezena de milhar
tmp(115)	:= "0101000000011";	-- STA @3                  	; armazena o novo valor do milhar
tmp(116)	:= "0110001011100";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(117)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(118)	:= "0101000000011";	-- STA @3                  	; armazena 0 no milhar
tmp(119)	:= "0001000000100";	-- LDA @4                  	; carrega o valor atual da dezena de milhar
tmp(120)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena de milhar
tmp(121)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(122)	:= "0111001111101";	-- JEQ .INCREMENTA_CMILHAR 	; se for, incrementa a centena de milhar
tmp(123)	:= "0101000000100";	-- STA @4                  	; armazena o novo valor da dezena de milhar
tmp(124)	:= "0110001011100";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(125)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(126)	:= "0101000000100";	-- STA @4                  	; armazena 0 na dezena de milhar
tmp(127)	:= "0001000000101";	-- LDA @5                  	; carrega o valor atual da centena de milhar
tmp(128)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena de milhar
tmp(129)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(130)	:= "0111010000101";	-- JEQ .INCREMENTA_MILHAO  	; se for, zera tudo
tmp(131)	:= "0101000000101";	-- STA @5                  	; armazena o novo valor da centena de milhar
tmp(132)	:= "0110001011100";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(133)	:= "0100000000000";	-- LDI $0  	; carrega 0
tmp(134)	:= "0101000000101";	-- STA $5  	; armazena 0 na centena de milhar
tmp(135)	:= "0110001011100";	-- JMP .FIM_INCREMENTA
tmp(136)	:= "0001000000000";	-- LDA @0      	; carrega o valor da unidade
tmp(137)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(138)	:= "0001000000001";	-- LDA @1      	; carrega o valor da dezena
tmp(139)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(140)	:= "0001000000010";	-- LDA @2      	; carrega o valor da centena
tmp(141)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(142)	:= "0001000000011";	-- LDA @3      	; carrega o valor do milhar
tmp(143)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(144)	:= "0001000000100";	-- LDA @4      	; carrega o valor da dezena de milhar
tmp(145)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(146)	:= "0001000000101";	-- LDA @5      	; carrega o valor da centena de milhar
tmp(147)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(148)	:= "1010000000000";	-- RET
tmp(149)	:= "0001000111001";	-- LDA @57                 	; carrega o intervalo atual
tmp(150)	:= "1000000001000";	-- CEQ @8                  	; verifica se é igual a 0
tmp(151)	:= "0111010100001";	-- JEQ .DIGITO_0_ML     	; se for
tmp(152)	:= "1000000001001";	-- CEQ @9                  	; verifica se é igual a 1
tmp(153)	:= "0111010101110";	-- JEQ .DIGITO_1_ML     	; se for
tmp(154)	:= "1000000001010";	-- CEQ @10                 	; verifica se é igual a 2
tmp(155)	:= "0111010111011";	-- JEQ .DIGITO_2_ML     	; se for
tmp(156)	:= "1000000001011";	-- CEQ @11                 	; verifica se é igual a 3
tmp(157)	:= "0111011001000";	-- JEQ .DIGITO_3_ML     	; se for
tmp(158)	:= "1000000001100";	-- CEQ @12                 	; verifica se é igual a 4
tmp(159)	:= "0111011010101";	-- JEQ .DIGITO_4_ML     	; se for
tmp(160)	:= "0110011100010";	-- JMP .DIGITO_5_ML 		; se não for nenhum dos acima
tmp(161)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(162)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(163)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(164)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(165)	:= "0001000111100";	-- LDA @60			; carrega o valor de centena do limite
tmp(166)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(167)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(168)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(169)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(170)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(171)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(172)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(173)	:= "1010000000000";	-- RET
tmp(174)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(175)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(176)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(177)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(178)	:= "0001000111100";	-- LDA @60     	; carrega o valor da centena do limite
tmp(179)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(180)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(181)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(182)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(183)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(184)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(185)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(186)	:= "1010000000000";	-- RET
tmp(187)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(188)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(189)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(190)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(191)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(192)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(193)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(194)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(195)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(196)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(197)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(198)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(199)	:= "1010000000000";	-- RET
tmp(200)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(201)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(202)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(203)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(204)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(205)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(206)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(207)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(208)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(209)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(210)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(211)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(212)	:= "1010000000000";	-- RET
tmp(213)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(214)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(215)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(216)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(217)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(218)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(219)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(220)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(221)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(222)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(223)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(224)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(225)	:= "1010000000000";	-- RET
tmp(226)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(227)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(228)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(229)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(230)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(231)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(232)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(233)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(234)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(235)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(236)	:= "0001101000000";	-- LDA @320     	; carrega o valor das chaves
tmp(237)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(238)	:= "1010000000000";	-- RET
tmp(239)	:= "0100000000000";	-- LDI $0
tmp(240)	:= "0101100000000";	-- STA @256
tmp(241)	:= "0101100000001";	-- STA @257
tmp(242)	:= "0101100000010";	-- STA @258
tmp(243)	:= "1010000000000";	-- RET
tmp(244)	:= "0001000111001";	-- LDA @57                 	; carrega o intervalo atual
tmp(245)	:= "1000000001000";	-- CEQ @8                  	; verifica se é igual a 0
tmp(246)	:= "0111100000000";	-- JEQ .DIGITO_0_MI     		; se for
tmp(247)	:= "1000000001001";	-- CEQ @9                  	; verifica se é igual a 1
tmp(248)	:= "0111100001010";	-- JEQ .DIGITO_1_MI     		; se for
tmp(249)	:= "1000000001010";	-- CEQ @10                 	; verifica se é igual a 2
tmp(250)	:= "0111100010100";	-- JEQ .DIGITO_2_MI     		; se for
tmp(251)	:= "1000000001011";	-- CEQ @11                 	; verifica se é igual a 3
tmp(252)	:= "0111100011110";	-- JEQ .DIGITO_3_MI     		; se for
tmp(253)	:= "1000000001100";	-- CEQ @12                 	; verifica se é igual a 4
tmp(254)	:= "0111100101001";	-- JEQ .DIGITO_4_MI     		; se for
tmp(255)	:= "0110100110011";	-- JMP .DIGITO_5_MI 			; se não for nenhum dos acima
tmp(256)	:= "0100000000001";	-- LDI $1			; atualiza o intervalo
tmp(257)	:= "0101000111001";	-- STA @57
tmp(258)	:= "0100000000110";	-- LDI $6			; acende os LEDs da segunda posição e apaga o resto
tmp(259)	:= "0101100000000";	-- STA @256
tmp(260)	:= "0100000000000";	-- LDI $0
tmp(261)	:= "0101100000001";	-- STA @257
tmp(262)	:= "0101100000010";	-- STA @258
tmp(263)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(264)	:= "0101000111010";	-- STA @58
tmp(265)	:= "1010000000000";	-- RET
tmp(266)	:= "0100000000010";	-- LDI $2			; atualiza o intervalo
tmp(267)	:= "0101000111001";	-- STA @57
tmp(268)	:= "0100000011000";	-- LDI $24			; acende os LEDs da terceira posição e apaga o resto
tmp(269)	:= "0101100000000";	-- STA @256
tmp(270)	:= "0100000000000";	-- LDI $0
tmp(271)	:= "0101100000001";	-- STA @257
tmp(272)	:= "0101100000010";	-- STA @258
tmp(273)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(274)	:= "0101000111011";	-- STA @59
tmp(275)	:= "1010000000000";	-- RET
tmp(276)	:= "0100000000011";	-- LDI $3			; atualiza o intervalo
tmp(277)	:= "0101000111001";	-- STA @57
tmp(278)	:= "0100001100000";	-- LDI $96			; acende os LEDs da quarta posição e apaga o resto
tmp(279)	:= "0101100000000";	-- STA @256
tmp(280)	:= "0100000000000";	-- LDI $0
tmp(281)	:= "0101100000001";	-- STA @257
tmp(282)	:= "0101100000010";	-- STA @258
tmp(283)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(284)	:= "0101000111100";	-- STA @60
tmp(285)	:= "1010000000000";	-- RET
tmp(286)	:= "0100000000100";	-- LDI $4			; atualiza o intervalo
tmp(287)	:= "0101000111001";	-- STA @57
tmp(288)	:= "0100010000000";	-- LDI $128		; acende os LEDs da quinta posição e apaga o resto
tmp(289)	:= "0101100000000";	-- STA @256
tmp(290)	:= "0100000000001";	-- LDI $1
tmp(291)	:= "0101100000001";	-- STA @257
tmp(292)	:= "0100000000000";	-- LDI $0
tmp(293)	:= "0101100000010";	-- STA @258
tmp(294)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(295)	:= "0101000111101";	-- STA @61
tmp(296)	:= "1010000000000";	-- RET
tmp(297)	:= "0100000000101";	-- LDI $5			; atualiza o intervalo
tmp(298)	:= "0101000111001";	-- STA @57
tmp(299)	:= "0100000000000";	-- LDI $0			; acende os LEDs da sexta posição e apaga o resto
tmp(300)	:= "0101100000000";	-- STA @256
tmp(301)	:= "0100000000001";	-- LDI $1
tmp(302)	:= "0101100000001";	-- STA @257
tmp(303)	:= "0101100000010";	-- STA @258
tmp(304)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(305)	:= "0101000111110";	-- STA @62
tmp(306)	:= "1010000000000";	-- RET
tmp(307)	:= "0100000000000";	-- LDI $0			; atualiza o intervalo
tmp(308)	:= "0101000111001";	-- STA @57
tmp(309)	:= "0100000000011";	-- LDI $3			; acende os LEDs da primeira posição e apaga o resto
tmp(310)	:= "0101100000000";	-- STA @256
tmp(311)	:= "0100000000000";	-- LDI $0
tmp(312)	:= "0101100000001";	-- STA @257
tmp(313)	:= "0101100000010";	-- STA @258
tmp(314)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(315)	:= "0101000111111";	-- STA @63
tmp(316)	:= "1010000000000";	-- RET
tmp(317)	:= "0001000000101";	-- LDA @5			; carrega o valor da centena de milhar
tmp(318)	:= "1000000111111";	-- CEQ @63			; compara com o valor limite da centena de milhar
tmp(319)	:= "0111101000010";	-- JEQ .CMILHAR_ATINGIU
tmp(320)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(321)	:= "1010000000000";	-- RET
tmp(322)	:= "0001000000100";	-- LDA @4			; carrega o valor da dezena de milhar
tmp(323)	:= "1000000111110";	-- CEQ @62			; compara com o valor limite da dezena de milhar
tmp(324)	:= "0111101000111";	-- JEQ .DMILHAR_ATINGIU
tmp(325)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(326)	:= "1010000000000";	-- RET
tmp(327)	:= "0001000000011";	-- LDA @3			; carrega o valor do milhar
tmp(328)	:= "1000000111101";	-- CEQ @61			; compara com o valor limite do milhar
tmp(329)	:= "0111101001100";	-- JEQ .MILHAR_ATINGIU
tmp(330)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(331)	:= "1010000000000";	-- RET
tmp(332)	:= "0001000000010";	-- LDA @2			; carrega o valor da centena
tmp(333)	:= "1000000111100";	-- CEQ @60			; compara com o valor limite da centena
tmp(334)	:= "0111101010001";	-- JEQ .CENTENA_ATINGIU
tmp(335)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(336)	:= "1010000000000";	-- RET
tmp(337)	:= "0001000000001";	-- LDA @1			; carrega o valor da dezena
tmp(338)	:= "1000000111011";	-- CEQ @59			; compara com o valor limite da dezena
tmp(339)	:= "0111101010110";	-- JEQ .DEZENA_ATINGIU
tmp(340)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(341)	:= "1010000000000";	-- RET
tmp(342)	:= "0001000000000";	-- LDA @0			; carrega o valor da unidade
tmp(343)	:= "1000000111010";	-- CEQ @58			; compara com o valor limite da unidade
tmp(344)	:= "0111101011011";	-- JEQ .UNIDADE_ATINGIU
tmp(345)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(346)	:= "1010000000000";	-- RET
tmp(347)	:= "0100000000001";	-- LDI $1
tmp(348)	:= "1010000000000";	-- RET
