tmp(0)	:= "0000000000000";	-- NOP
tmp(1)	:= "0001000000000";	-- LDA $0
tmp(2)	:= "0101100100000";	-- STA @288
tmp(3)	:= "0010000000001";	-- ADD $1
tmp(4)	:= "0110000000101";	-- JMP .TEST
tmp(5)	:= "0110000000110";	-- JMP .TEST2
tmp(6)	:= "0110000000000";	-- JMP .LOOP
