tmp(0)	:= "0000000000000";	-- 	; SETUP
tmp(1)	:= "0101111111111";	-- STA @511    	; reseta a leitura do key 0
tmp(2)	:= "0101111111110";	-- STA @510    	; reseta a leitura do key 1
tmp(3)	:= "0101111111101";	-- STA @509    	; reseta a leitura do key reset
tmp(4)	:= "0100000000000";	-- LDI $0      	; carrega o valor inicial das casas
tmp(5)	:= "0101000111001";	-- STA @57     	; intervalo numérico de configuração
tmp(6)	:= "0101000000000";	-- STA @0      	; armazena 0 na unidade
tmp(7)	:= "0101000000001";	-- STA @1      	; armazena 0 na dezena
tmp(8)	:= "0101000000010";	-- STA @2      	; armazena 0 na centena
tmp(9)	:= "0101000000011";	-- STA @3      	; armazena 0 no milhar
tmp(10)	:= "0101000000100";	-- STA @4      	; armazena 0 na dezena de milhar
tmp(11)	:= "0101000000101";	-- STA @5      	; armazena 0 na centena de milhar
tmp(12)	:= "0101000001000";	-- STA @8      	; armazena um 0 de referência
tmp(13)	:= "0100000000001";	-- LDI $1      	; carrega o valor de incremento
tmp(14)	:= "0101000000110";	-- STA @6      	; armazena o valor de incremento
tmp(15)	:= "0101000001001";	-- STA @9			; armazena 1 no 9 para referência do intervalo numérico de configuração
tmp(16)	:= "0100000001010";	-- LDI $10     	; carrega o valor máximo por casa possível
tmp(17)	:= "0101000000111";	-- STA @7      	; armazena o valor máximo por casa possível
tmp(18)	:= "0100000001001";	-- LDI $9      	; carrega o número 9 para definir o limite de contagem inicial
tmp(19)	:= "0101000111010";	-- STA @58     	; armazena na casa das unidades do limite
tmp(20)	:= "0101000111011";	-- STA @59     	; armazena na casa das dezenas do limite
tmp(21)	:= "0101000111100";	-- STA @60     	; armazena na casa das centenas do limite
tmp(22)	:= "0101000111101";	-- STA @61     	; armazena na casa dos milhares do limite
tmp(23)	:= "0101000111110";	-- STA @62     	; armazena na casa das dezenas de milhar do limite
tmp(24)	:= "0101000111111";	-- STA @63     	; armazena na casa das centenas de milhar do limite
tmp(25)	:= "0100000000010";	-- LDI $2			; carrega 2 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(26)	:= "0101000001010";	-- STA @10			; armazena a referência de estado 2 no endereço 10
tmp(27)	:= "0100000000011";	-- LDI $3			; carrega 3 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(28)	:= "0101000001011";	-- STA @11			; armazena a referência de estado 3 no endereço 11
tmp(29)	:= "0100000000100";	-- LDI $4			; carrega 4 para inicializar próximo endereço de referência do intervalo numérico de configuração
tmp(30)	:= "0101000001100";	-- STA @12			; armazena a referência de estado 4 no endereço 12
tmp(31)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(32)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(33)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(34)	:= "0111000100101";	-- JEQ .PULA_RESET
tmp(35)	:= "0101111111101";	-- STA @509
tmp(36)	:= "1001001010010";	-- JSR .RESET
tmp(37)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(38)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(39)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(40)	:= "0111000101011";	-- JEQ .PULA_CONFIG
tmp(41)	:= "0101111111110";	-- STA @510
tmp(42)	:= "0110000110110";	-- JMP .INICIO_LOOP_CONFIGURACAO_LIMITE
tmp(43)	:= "1001101000111";	-- JSR .ATINGIU_LIMITE			; verifica se a contagem atingiu o limite
tmp(44)	:= "1000000000110";	-- CEQ @6						; se atingiu o limite, pula o incrementa contagem
tmp(45)	:= "0111000110100";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(46)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(47)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(48)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(49)	:= "0111000110100";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(50)	:= "0101111111111";	-- STA @511
tmp(51)	:= "1001001100001";	-- JSR .INCREMENTA_CONTAGEM
tmp(52)	:= "1001010010010";	-- JSR .MOSTRA_CONTAGEM    	; escreve os números da contagem nos displays
tmp(53)	:= "0110000011111";	-- JMP .LOOP_PRINCIPAL
tmp(54)	:= "1001001010010";	-- JSR .RESET		; reseta a contagem
tmp(55)	:= "0100000000011";	-- LDI $3			; acende os leds da primeira posição
tmp(56)	:= "0101100000000";	-- STA @256
tmp(57)	:= "0100000000000";	-- LDI $0
tmp(58)	:= "0101100000001";	-- STA @257
tmp(59)	:= "0101100000010";	-- STA @258
tmp(60)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(61)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(62)	:= "1000000000110";	-- CEQ @6      	; verifica se é 1
tmp(63)	:= "0111001001110";	-- JEQ .SAIR_LOOP_CONFIGURACAO_LIMITE
tmp(64)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(65)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(66)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(67)	:= "0111001000110";	-- JEQ .PULA_MUDANCA_ESTADO
tmp(68)	:= "0101111111110";	-- STA @510
tmp(69)	:= "0110001001110";	-- JMP .SAIR_LOOP_CONFIGURACAO_LIMITE
tmp(70)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(71)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(72)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(73)	:= "0111001001100";	-- JEQ .PULA_MUDANCA_INTERVALO
tmp(74)	:= "0101111111111";	-- STA @511
tmp(75)	:= "1001011111110";	-- JSR .MUDA_INTERVALO
tmp(76)	:= "1001010011111";	-- JSR .MOSTRA_LIMITE
tmp(77)	:= "0110000111100";	-- JMP .LOOP_CONFIGURACAO_LIMITE
tmp(78)	:= "1001011111001";	-- JSR .APAGA_LEDS         	; apaga os LEDs
tmp(79)	:= "0100000000000";	-- LDI $0    		; carrega 0
tmp(80)	:= "0101000111001";	-- STA @57     	; armazena 0 no intervalo de mudança atual
tmp(81)	:= "0110000011111";	-- JMP .LOOP_PRINCIPAL
tmp(82)	:= "0100000000000";	-- LDI $0
tmp(83)	:= "0101000000000";	-- STA @0
tmp(84)	:= "0101000000001";	-- STA @1
tmp(85)	:= "0101000000010";	-- STA @2
tmp(86)	:= "0101000000011";	-- STA @3
tmp(87)	:= "0101000000100";	-- STA @4
tmp(88)	:= "0101000000101";	-- STA @5
tmp(89)	:= "0100000000000";	-- LDI $0
tmp(90)	:= "0101100000000";	-- STA @256
tmp(91)	:= "0101100000001";	-- STA @257
tmp(92)	:= "0101100000010";	-- STA @258
tmp(93)	:= "0101111111111";	-- STA @511
tmp(94)	:= "0101111111110";	-- STA @510
tmp(95)	:= "0101111111101";	-- STA @509
tmp(96)	:= "1010000000000";	-- RET
tmp(97)	:= "0001000000000";	-- LDA @0                  	; carrega o valor da unidade
tmp(98)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da unidade
tmp(99)	:= "1000000000111";	-- CEQ @7                  	; compara o valor da casa com 10
tmp(100)	:= "0111001100111";	-- JEQ .INCREMENTA_DEZENA  	; incrementa a casa da dezena caso necessário
tmp(101)	:= "0101000000000";	-- STA @0                  	; armazena o valor da unidade
tmp(102)	:= "1010000000000";	-- RET
tmp(103)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(104)	:= "0101000000000";	-- STA @0                  	; armazena 0 na unidade
tmp(105)	:= "0001000000001";	-- LDA @1                  	; carrega o valor atual da dezena
tmp(106)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena
tmp(107)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(108)	:= "0111001101111";	-- JEQ .INCREMENTA_CENTENA 	; se for, incrementa a centena
tmp(109)	:= "0101000000001";	-- STA @1                  	; armazena o novo valor da dezena
tmp(110)	:= "0110001100110";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(111)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(112)	:= "0101000000001";	-- STA @1                  	; armazena 0 na dezena
tmp(113)	:= "0001000000010";	-- LDA @2                  	; carrega o valor atual da centena
tmp(114)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena
tmp(115)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(116)	:= "0111001110111";	-- JEQ .INCREMENTA_MILHAR  	; se for, incrementa o milhar
tmp(117)	:= "0101000000010";	-- STA @2                  	; armazena o novo valor da centena
tmp(118)	:= "0110001100110";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(119)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(120)	:= "0101000000010";	-- STA @2                  	; armazena 0 na centena
tmp(121)	:= "0001000000011";	-- LDA @3                  	; carrega o valor atual do milhar
tmp(122)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor do milhar
tmp(123)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(124)	:= "0111001111111";	-- JEQ .INCREMENTA_DMILHAR 	; se for, incrementa a dezena de milhar
tmp(125)	:= "0101000000011";	-- STA @3                  	; armazena o novo valor do milhar
tmp(126)	:= "0110001100110";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(127)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(128)	:= "0101000000011";	-- STA @3                  	; armazena 0 no milhar
tmp(129)	:= "0001000000100";	-- LDA @4                  	; carrega o valor atual da dezena de milhar
tmp(130)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena de milhar
tmp(131)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(132)	:= "0111010000111";	-- JEQ .INCREMENTA_CMILHAR 	; se for, incrementa a centena de milhar
tmp(133)	:= "0101000000100";	-- STA @4                  	; armazena o novo valor da dezena de milhar
tmp(134)	:= "0110001100110";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(135)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(136)	:= "0101000000100";	-- STA @4                  	; armazena 0 na dezena de milhar
tmp(137)	:= "0001000000101";	-- LDA @5                  	; carrega o valor atual da centena de milhar
tmp(138)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena de milhar
tmp(139)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(140)	:= "0111010001111";	-- JEQ .INCREMENTA_MILHAO  	; se for, zera tudo
tmp(141)	:= "0101000000101";	-- STA @5                  	; armazena o novo valor da centena de milhar
tmp(142)	:= "0110001100110";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(143)	:= "0100000000000";	-- LDI $0  	; carrega 0
tmp(144)	:= "0101000000101";	-- STA $5  	; armazena 0 na centena de milhar
tmp(145)	:= "0110001100110";	-- JMP .FIM_INCREMENTA
tmp(146)	:= "0001000000000";	-- LDA @0      	; carrega o valor da unidade
tmp(147)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(148)	:= "0001000000001";	-- LDA @1      	; carrega o valor da dezena
tmp(149)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(150)	:= "0001000000010";	-- LDA @2      	; carrega o valor da centena
tmp(151)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(152)	:= "0001000000011";	-- LDA @3      	; carrega o valor do milhar
tmp(153)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(154)	:= "0001000000100";	-- LDA @4      	; carrega o valor da dezena de milhar
tmp(155)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(156)	:= "0001000000101";	-- LDA @5      	; carrega o valor da centena de milhar
tmp(157)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(158)	:= "1010000000000";	-- RET
tmp(159)	:= "0001000111001";	-- LDA @57                 	; carrega o intervalo atual
tmp(160)	:= "1000000001000";	-- CEQ @8                  	; verifica se é igual a 0
tmp(161)	:= "0111010101011";	-- JEQ .DIGITO_0_ML     	; se for
tmp(162)	:= "1000000001001";	-- CEQ @9                  	; verifica se é igual a 1
tmp(163)	:= "0111010111000";	-- JEQ .DIGITO_1_ML     	; se for
tmp(164)	:= "1000000001010";	-- CEQ @10                 	; verifica se é igual a 2
tmp(165)	:= "0111011000101";	-- JEQ .DIGITO_2_ML     	; se for
tmp(166)	:= "1000000001011";	-- CEQ @11                 	; verifica se é igual a 3
tmp(167)	:= "0111011010010";	-- JEQ .DIGITO_3_ML     	; se for
tmp(168)	:= "1000000001100";	-- CEQ @12                 	; verifica se é igual a 4
tmp(169)	:= "0111011011111";	-- JEQ .DIGITO_4_ML     	; se for
tmp(170)	:= "0110011101100";	-- JMP .DIGITO_5_ML 		; se não for nenhum dos acima
tmp(171)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(172)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(173)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(174)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(175)	:= "0001000111100";	-- LDA @60			; carrega o valor de centena do limite
tmp(176)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(177)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(178)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(179)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(180)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(181)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(182)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(183)	:= "1010000000000";	-- RET
tmp(184)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(185)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(186)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(187)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(188)	:= "0001000111100";	-- LDA @60     	; carrega o valor da centena do limite
tmp(189)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(190)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(191)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(192)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(193)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(194)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(195)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(196)	:= "1010000000000";	-- RET
tmp(197)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(198)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(199)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(200)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(201)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(202)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(203)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(204)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(205)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(206)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(207)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(208)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(209)	:= "1010000000000";	-- RET
tmp(210)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(211)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(212)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(213)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(214)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(215)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(216)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(217)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(218)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(219)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(220)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(221)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(222)	:= "1010000000000";	-- RET
tmp(223)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(224)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(225)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(226)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(227)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(228)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(229)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(230)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(231)	:= "0001101000000";	-- LDA @320    	; carrega o valor das chaves
tmp(232)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(233)	:= "0001000111111";	-- LDA @63     	; carrega o valor da centena de milhar do limite
tmp(234)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(235)	:= "1010000000000";	-- RET
tmp(236)	:= "0001000111010";	-- LDA @58     	; carrega o valor da unidade do limite
tmp(237)	:= "0101100100000";	-- STA @288    	; armazena no HEX 0
tmp(238)	:= "0001000111011";	-- LDA @59			; carrega o valor da dezena do limite
tmp(239)	:= "0101100100001";	-- STA @289    	; armazena no HEX 1
tmp(240)	:= "0001000111100";	-- LDA @60    		; carrega o valor da centena do limite
tmp(241)	:= "0101100100010";	-- STA @290    	; armazena no HEX 2
tmp(242)	:= "0001000111101";	-- LDA @61     	; carrega o valor do milhar do limite
tmp(243)	:= "0101100100011";	-- STA @291    	; armazena no HEX 3
tmp(244)	:= "0001000111110";	-- LDA @62     	; carrega o valor da dezena de milhar do limite
tmp(245)	:= "0101100100100";	-- STA @292    	; armazena no HEX 4
tmp(246)	:= "0001101000000";	-- LDA @320     	; carrega o valor das chaves
tmp(247)	:= "0101100100101";	-- STA @293    	; armazena no HEX 5
tmp(248)	:= "1010000000000";	-- RET
tmp(249)	:= "0100000000000";	-- LDI $0
tmp(250)	:= "0101100000000";	-- STA @256
tmp(251)	:= "0101100000001";	-- STA @257
tmp(252)	:= "0101100000010";	-- STA @258
tmp(253)	:= "1010000000000";	-- RET
tmp(254)	:= "0001000111001";	-- LDA @57                 	; carrega o intervalo atual
tmp(255)	:= "1000000001000";	-- CEQ @8                  	; verifica se é igual a 0
tmp(256)	:= "0111100001010";	-- JEQ .DIGITO_0_MI     		; se for
tmp(257)	:= "1000000001001";	-- CEQ @9                  	; verifica se é igual a 1
tmp(258)	:= "0111100010100";	-- JEQ .DIGITO_1_MI     		; se for
tmp(259)	:= "1000000001010";	-- CEQ @10                 	; verifica se é igual a 2
tmp(260)	:= "0111100011110";	-- JEQ .DIGITO_2_MI     		; se for
tmp(261)	:= "1000000001011";	-- CEQ @11                 	; verifica se é igual a 3
tmp(262)	:= "0111100101000";	-- JEQ .DIGITO_3_MI     		; se for
tmp(263)	:= "1000000001100";	-- CEQ @12                 	; verifica se é igual a 4
tmp(264)	:= "0111100110011";	-- JEQ .DIGITO_4_MI     		; se for
tmp(265)	:= "0110100111101";	-- JMP .DIGITO_5_MI 			; se não for nenhum dos acima
tmp(266)	:= "0100000000001";	-- LDI $1			; atualiza o intervalo
tmp(267)	:= "0101000111001";	-- STA @57
tmp(268)	:= "0100000000110";	-- LDI $6			; acende os LEDs da segunda posição e apaga o resto
tmp(269)	:= "0101100000000";	-- STA @256
tmp(270)	:= "0100000000000";	-- LDI $0
tmp(271)	:= "0101100000001";	-- STA @257
tmp(272)	:= "0101100000010";	-- STA @258
tmp(273)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(274)	:= "0101000111010";	-- STA @58
tmp(275)	:= "1010000000000";	-- RET
tmp(276)	:= "0100000000010";	-- LDI $2			; atualiza o intervalo
tmp(277)	:= "0101000111001";	-- STA @57
tmp(278)	:= "0100000011000";	-- LDI $24			; acende os LEDs da terceira posição e apaga o resto
tmp(279)	:= "0101100000000";	-- STA @256
tmp(280)	:= "0100000000000";	-- LDI $0
tmp(281)	:= "0101100000001";	-- STA @257
tmp(282)	:= "0101100000010";	-- STA @258
tmp(283)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(284)	:= "0101000111011";	-- STA @59
tmp(285)	:= "1010000000000";	-- RET
tmp(286)	:= "0100000000011";	-- LDI $3			; atualiza o intervalo
tmp(287)	:= "0101000111001";	-- STA @57
tmp(288)	:= "0100001100000";	-- LDI $96			; acende os LEDs da quarta posição e apaga o resto
tmp(289)	:= "0101100000000";	-- STA @256
tmp(290)	:= "0100000000000";	-- LDI $0
tmp(291)	:= "0101100000001";	-- STA @257
tmp(292)	:= "0101100000010";	-- STA @258
tmp(293)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(294)	:= "0101000111100";	-- STA @60
tmp(295)	:= "1010000000000";	-- RET
tmp(296)	:= "0100000000100";	-- LDI $4			; atualiza o intervalo
tmp(297)	:= "0101000111001";	-- STA @57
tmp(298)	:= "0100010000000";	-- LDI $128		; acende os LEDs da quinta posição e apaga o resto
tmp(299)	:= "0101100000000";	-- STA @256
tmp(300)	:= "0100000000001";	-- LDI $1
tmp(301)	:= "0101100000001";	-- STA @257
tmp(302)	:= "0100000000000";	-- LDI $0
tmp(303)	:= "0101100000010";	-- STA @258
tmp(304)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(305)	:= "0101000111101";	-- STA @61
tmp(306)	:= "1010000000000";	-- RET
tmp(307)	:= "0100000000101";	-- LDI $5			; atualiza o intervalo
tmp(308)	:= "0101000111001";	-- STA @57
tmp(309)	:= "0100000000000";	-- LDI $0			; acende os LEDs da sexta posição e apaga o resto
tmp(310)	:= "0101100000000";	-- STA @256
tmp(311)	:= "0100000000001";	-- LDI $1
tmp(312)	:= "0101100000001";	-- STA @257
tmp(313)	:= "0101100000010";	-- STA @258
tmp(314)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(315)	:= "0101000111110";	-- STA @62
tmp(316)	:= "1010000000000";	-- RET
tmp(317)	:= "0100000000000";	-- LDI $0			; atualiza o intervalo
tmp(318)	:= "0101000111001";	-- STA @57
tmp(319)	:= "0100000000011";	-- LDI $3			; acende os LEDs da primeira posição e apaga o resto
tmp(320)	:= "0101100000000";	-- STA @256
tmp(321)	:= "0100000000000";	-- LDI $0
tmp(322)	:= "0101100000001";	-- STA @257
tmp(323)	:= "0101100000010";	-- STA @258
tmp(324)	:= "0001101000000";	-- LDA @320		; salva o novo valor do dígito
tmp(325)	:= "0101000111111";	-- STA @63
tmp(326)	:= "1010000000000";	-- RET
tmp(327)	:= "0001000000101";	-- LDA @5			; carrega o valor da centena de milhar
tmp(328)	:= "1000000111111";	-- CEQ @63			; compara com o valor limite da centena de milhar
tmp(329)	:= "0111101001100";	-- JEQ .CMILHAR_ATINGIU
tmp(330)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(331)	:= "1010000000000";	-- RET
tmp(332)	:= "0001000000100";	-- LDA @4			; carrega o valor da dezena de milhar
tmp(333)	:= "1000000111110";	-- CEQ @62			; compara com o valor limite da dezena de milhar
tmp(334)	:= "0111101010001";	-- JEQ .DMILHAR_ATINGIU
tmp(335)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(336)	:= "1010000000000";	-- RET
tmp(337)	:= "0001000000011";	-- LDA @3			; carrega o valor do milhar
tmp(338)	:= "1000000111101";	-- CEQ @61			; compara com o valor limite do milhar
tmp(339)	:= "0111101010110";	-- JEQ .MILHAR_ATINGIU
tmp(340)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(341)	:= "1010000000000";	-- RET
tmp(342)	:= "0001000000010";	-- LDA @2			; carrega o valor da centena
tmp(343)	:= "1000000111100";	-- CEQ @60			; compara com o valor limite da centena
tmp(344)	:= "0111101011011";	-- JEQ .CENTENA_ATINGIU
tmp(345)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(346)	:= "1010000000000";	-- RET
tmp(347)	:= "0001000000001";	-- LDA @1			; carrega o valor da dezena
tmp(348)	:= "1000000111011";	-- CEQ @59			; compara com o valor limite da dezena
tmp(349)	:= "0111101100000";	-- JEQ .DEZENA_ATINGIU
tmp(350)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(351)	:= "1010000000000";	-- RET
tmp(352)	:= "0001000000000";	-- LDA @0			; carrega o valor da unidade
tmp(353)	:= "1000000111010";	-- CEQ @58			; compara com o valor limite da unidade
tmp(354)	:= "0111101100101";	-- JEQ .UNIDADE_ATINGIU
tmp(355)	:= "0100000000000";	-- LDI $0			; se não for igual, não atingiu
tmp(356)	:= "1010000000000";	-- RET
tmp(357)	:= "0100011111111";	-- LDI $255
tmp(358)	:= "0101100000000";	-- STA @256
tmp(359)	:= "0101100000001";	-- STA @257
tmp(360)	:= "0101100000010";	-- STA @258
tmp(361)	:= "0100000000001";	-- LDI $1
tmp(362)	:= "1010000000000";	-- RET
