tmp(0)	:= "0000000000000";	-- 	; SETUP
tmp(1)	:= "0000000000000";	-- NOP
tmp(2)	:= "0101111111111";	-- STA @511    	; reseta a leitura do key 0
tmp(3)	:= "0101111111110";	-- STA @510    	; reseta a leitura do key 1
tmp(4)	:= "0101111111101";	-- STA @509    	; reseta a leitura do key reset
tmp(5)	:= "0100000000000";	-- LDI $0      	; carrega o valor inicial das casas
tmp(6)	:= "0101000000000";	-- STA @0      	; armazena 0 na unidade
tmp(7)	:= "0101000000001";	-- STA @1      	; armazena 0 na dezena
tmp(8)	:= "0101000000010";	-- STA @2      	; armazena 0 na centena
tmp(9)	:= "0101000000011";	-- STA @3      	; armazena 0 no milhar
tmp(10)	:= "0101000000100";	-- STA @4      	; armazena 0 na dezena de milhar
tmp(11)	:= "0101000000101";	-- STA @5      	; armazena 0 na centena de milhar
tmp(12)	:= "0101000001000";	-- STA @8      	; armazena um 0 de referência
tmp(13)	:= "0100000000001";	-- LDI $1      	; carrega o valor de incremento
tmp(14)	:= "0101000000110";	-- STA @6      	; armazena o valor de incremento
tmp(15)	:= "0100000001010";	-- LDI $10     	; carrega o valor máximo por casa possível
tmp(16)	:= "0101000000111";	-- STA @7      	; armazena o valor máximo por casa possível
tmp(17)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(18)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(19)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(20)	:= "0111000010111";	-- JEQ .PULA_RESET
tmp(21)	:= "0101111111101";	-- STA @509
tmp(22)	:= "1001000110110";	-- JSR .RESET
tmp(23)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(24)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(25)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(26)	:= "0111000011101";	-- JEQ .PULA_CONFIG
tmp(27)	:= "0101111111110";	-- STA @510
tmp(28)	:= "0110000100111";	-- JMP .LOOP_CONFIGURACAO_LIMITE
tmp(29)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(30)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(31)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(32)	:= "0111000100011";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(33)	:= "0101111111111";	-- STA @511
tmp(34)	:= "1001000111110";	-- JSR .INCREMENTA_CONTAGEM
tmp(35)	:= "0100000000000";	-- LDI $0                  	; define se apaga ou acende os LEDS
tmp(36)	:= "1001001111100";	-- JSR .MODIFICA_LEDS      	; apaga os LEDs
tmp(37)	:= "1001001101111";	-- JSR .MOSTRA_CONTAGEM    	; escreve os números da contagem nos displays
tmp(38)	:= "0110000010001";	-- JMP .LOOP_PRINCIPAL
tmp(39)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(40)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(41)	:= "1000000000110";	-- CEQ @6      	; verifica se é 1
tmp(42)	:= "0111000010001";	-- JEQ .LOOP_PRINCIPAL
tmp(43)	:= "0001101100001";	-- LDA @353    	; carrega o valor do botão 1
tmp(44)	:= "1011000000110";	-- AND @6      	; aplica a mask
tmp(45)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(46)	:= "0111000110010";	-- JEQ .PULA_MUDANCA
tmp(47)	:= "0101111111110";	-- STA @510
tmp(48)	:= "0101111111111";	-- STA @511
tmp(49)	:= "0110000010001";	-- JMP .LOOP_PRINCIPAL
tmp(50)	:= "0100011111111";	-- LDI $255
tmp(51)	:= "1001001111100";	-- JSR .MODIFICA_LEDS
tmp(52)	:= "0110000100111";	-- JMP .LOOP_CONFIGURACAO_LIMITE
tmp(53)	:= "0110000110101";	-- JMP .FIM
tmp(54)	:= "0100000000000";	-- LDI $0
tmp(55)	:= "0101000000000";	-- STA @0
tmp(56)	:= "0101000000001";	-- STA @1
tmp(57)	:= "0101000000010";	-- STA @2
tmp(58)	:= "0101000000011";	-- STA @3
tmp(59)	:= "0101000000100";	-- STA @4
tmp(60)	:= "0101000000101";	-- STA @5
tmp(61)	:= "1000000000000";	-- RET
tmp(62)	:= "0001000000000";	-- LDA @0                  	; carrega o valor da unidade
tmp(63)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da unidade
tmp(64)	:= "1000000000111";	-- CEQ @7                  	; compara o valor da casa com 10
tmp(65)	:= "0111001000100";	-- JEQ .INCREMENTA_DEZENA  	; incrementa a casa da dezena caso necessário
tmp(66)	:= "0101000000000";	-- STA @0                  	; armazena o valor da unidade
tmp(67)	:= "1000000000000";	-- RET
tmp(68)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(69)	:= "0101000000000";	-- STA @0                  	; armazena 0 na unidade
tmp(70)	:= "0001000000001";	-- LDA @1                  	; carrega o valor atual da dezena
tmp(71)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena
tmp(72)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(73)	:= "0111001001100";	-- JEQ .INCREMENTA_CENTENA 	; se for, incrementa a centena
tmp(74)	:= "0101000000001";	-- STA @1                  	; armazena o novo valor da dezena
tmp(75)	:= "0110001000011";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(76)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(77)	:= "0101000000001";	-- STA @1                  	; armazena 0 na dezena
tmp(78)	:= "0001000000010";	-- LDA @2                  	; carrega o valor atual da centena
tmp(79)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena
tmp(80)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(81)	:= "0111001010100";	-- JEQ .INCREMENTA_MILHAR  	; se for, incrementa o milhar
tmp(82)	:= "0101000000010";	-- STA @2                  	; armazena o novo valor da centena
tmp(83)	:= "0110001000011";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(84)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(85)	:= "0101000000010";	-- STA @2                  	; armazena 0 na centena
tmp(86)	:= "0001000000011";	-- LDA @3                  	; carrega o valor atual do milhar
tmp(87)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor do milhar
tmp(88)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(89)	:= "0111001011100";	-- JEQ .INCREMENTA_DMILHAR 	; se for, incrementa a dezena de milhar
tmp(90)	:= "0101000000011";	-- STA @3                  	; armazena o novo valor do milhar
tmp(91)	:= "0110001000011";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(92)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(93)	:= "0101000000011";	-- STA @3                  	; armazena 0 no milhar
tmp(94)	:= "0001000000100";	-- LDA @4                  	; carrega o valor atual da dezena de milhar
tmp(95)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena de milhar
tmp(96)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(97)	:= "0111001100100";	-- JEQ .INCREMENTA_CMILHAR 	; se for, incrementa a centena de milhar
tmp(98)	:= "0101000000100";	-- STA @4                  	; armazena o novo valor da dezena de milhar
tmp(99)	:= "0110001000011";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(100)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(101)	:= "0101000000100";	-- STA @4                  	; armazena 0 na dezena de milhar
tmp(102)	:= "0001000000101";	-- LDA @5                  	; carrega o valor atual da centena de milhar
tmp(103)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena de milhar
tmp(104)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(105)	:= "0111001101100";	-- JEQ .INCREMENTA_MILHAO  	; se for, zera tudo
tmp(106)	:= "0101000000101";	-- STA @5                  	; armazena o novo valor da centena de milhar
tmp(107)	:= "0110001000011";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(108)	:= "0100000000000";	-- LDI $0  	; carrega 0
tmp(109)	:= "0101000000101";	-- STA $5  	; armazena 0 na centena de milhar
tmp(110)	:= "0110001000011";	-- JMP .FIM_INCREMENTA
tmp(111)	:= "0001000000000";	-- LDA @0      	; carrega o valor da unidade
tmp(112)	:= "0101100100000";	-- STA @288    	; armazena o 0 no HEX 0
tmp(113)	:= "0001000000001";	-- LDA @1      	; carrega o valor da dezena
tmp(114)	:= "0101100100001";	-- STA @289    	; armazena o 0 no HEX 1
tmp(115)	:= "0001000000010";	-- LDA @2      	; carrega o valor da centena
tmp(116)	:= "0101100100010";	-- STA @290    	; armazena o 0 no HEX 2
tmp(117)	:= "0001000000011";	-- LDA @3      	; carrega o valor do milhar
tmp(118)	:= "0101100100011";	-- STA @291    	; armazena o 0 no HEX 3
tmp(119)	:= "0001000000100";	-- LDA @4      	; carrega o valor da dezena de milhar
tmp(120)	:= "0101100100100";	-- STA @292    	; armazena o 0 no HEX 4
tmp(121)	:= "0001000000101";	-- LDA @5      	; carrega o valor da centena de milhar
tmp(122)	:= "0101100100101";	-- STA @293    	; armazena o 0 no HEX 5
tmp(123)	:= "1000000000000";	-- RET
tmp(124)	:= "0101100000000";	-- STA @256
tmp(125)	:= "0101100000001";	-- STA @257
tmp(126)	:= "0101100000010";	-- STA @258
tmp(127)	:= "1000000000000";	-- RET
