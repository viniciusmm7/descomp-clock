tmp(0)	:= "0000000000000";	-- 	; SETUP
tmp(1)	:= "0000000000000";	-- NOP
tmp(2)	:= "0101111111111";	-- STA @511    	; reseta a leitura do key 0
tmp(3)	:= "0101111111110";	-- STA @510    	; reseta a leitura do key 1
tmp(4)	:= "0101111111101";	-- STA @509    	; reseta a leitura do key reset
tmp(5)	:= "0100000000000";	-- LDI $0      	; carrega o valor inicial das casas
tmp(6)	:= "0101000000000";	-- STA @0      	; armazena 0 na unidade
tmp(7)	:= "0101000000001";	-- STA @1      	; armazena 0 na dezena
tmp(8)	:= "0101000000010";	-- STA @2      	; armazena 0 na centena
tmp(9)	:= "0101000000011";	-- STA @3      	; armazena 0 no milhar
tmp(10)	:= "0101000000100";	-- STA @4      	; armazena 0 na dezena de milhar
tmp(11)	:= "0101000000101";	-- STA @5      	; armazena 0 na centena de milhar
tmp(12)	:= "0101000001000";	-- STA @8      	; armazena um 0 de referência
tmp(13)	:= "0100000000001";	-- LDI $1      	; carrega o valor de incremento
tmp(14)	:= "0101000000110";	-- STA @6      	; armazena o valor de incremento
tmp(15)	:= "0100000001010";	-- LDI $10     	; carrega o valor máximo por casa possível
tmp(16)	:= "0101000000111";	-- STA @7      	; armazena o valor máximo por casa possível
tmp(17)	:= "0001101100100";	-- LDA @356    	; carrega o valor do botão reset
tmp(18)	:= "11@6000000000";	-- AND @6      	; aplica a mask
tmp(19)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(20)	:= "0111000010111";	-- JEQ .PULA_RESET
tmp(21)	:= "0101111111101";	-- STA @509
tmp(22)	:= "1001000100000";	-- JSR .RESET
tmp(23)	:= "0001101100000";	-- LDA @352    	; carrega o valor do botão 0
tmp(24)	:= "11@6000000000";	-- AND @6      	; aplica a mask
tmp(25)	:= "1000000001000";	-- CEQ @8      	; verifica se é 0
tmp(26)	:= "0111000011101";	-- JEQ .PULA_INCREMENTA_CONTAGEM
tmp(27)	:= "0101111111111";	-- STA @511
tmp(28)	:= "1001000101000";	-- JSR .INCREMENTA_CONTAGEM
tmp(29)	:= "1001001011001";	-- JSR .ATUALIZA_DISPLAYS
tmp(30)	:= "0110000010001";	-- JMP .LOOP
tmp(31)	:= "0110000011111";	-- JMP .FIM
tmp(32)	:= "0100000000000";	-- LDI $0
tmp(33)	:= "0101000000000";	-- STA @0
tmp(34)	:= "0101000000001";	-- STA @1
tmp(35)	:= "0101000000010";	-- STA @2
tmp(36)	:= "0101000000011";	-- STA @3
tmp(37)	:= "0101000000100";	-- STA @4
tmp(38)	:= "0101000000101";	-- STA @5
tmp(39)	:= "1000000000000";	-- RET
tmp(40)	:= "0001000000000";	-- LDA @0                  	; carrega o valor da unidade
tmp(41)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da unidade
tmp(42)	:= "1000000000111";	-- CEQ @7                  	; compara o valor da casa com 10
tmp(43)	:= "0111000101110";	-- JEQ .INCREMENTA_DEZENA  	; incrementa a casa da dezena caso necessário
tmp(44)	:= "0101000000000";	-- STA @0                  	; armazena o valor da unidade
tmp(45)	:= "1000000000000";	-- RET
tmp(46)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(47)	:= "0101000000000";	-- STA @0                  	; armazena 0 na unidade
tmp(48)	:= "0001000000001";	-- LDA @1                  	; carrega o valor atual da dezena
tmp(49)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena
tmp(50)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(51)	:= "0111000110110";	-- JEQ .INCREMENTA_CENTENA 	; se for, incrementa a centena
tmp(52)	:= "0101000000001";	-- STA @1                  	; armazena o novo valor da dezena
tmp(53)	:= "0110000101101";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(54)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(55)	:= "0101000000001";	-- STA @1                  	; armazena 0 na dezena
tmp(56)	:= "0001000000010";	-- LDA @2                  	; carrega o valor atual da centena
tmp(57)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena
tmp(58)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(59)	:= "0111000111110";	-- JEQ .INCREMENTA_MILHAR  	; se for, incrementa o milhar
tmp(60)	:= "0101000000010";	-- STA @2                  	; armazena o novo valor da centena
tmp(61)	:= "0110000101101";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(62)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(63)	:= "0101000000010";	-- STA @2                  	; armazena 0 na centena
tmp(64)	:= "0001000000011";	-- LDA @3                  	; carrega o valor atual do milhar
tmp(65)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor do milhar
tmp(66)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(67)	:= "0111001000110";	-- JEQ .INCREMENTA_DMILHAR 	; se for, incrementa a dezena de milhar
tmp(68)	:= "0101000000011";	-- STA @3                  	; armazena o novo valor do milhar
tmp(69)	:= "0110000101101";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(70)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(71)	:= "0101000000011";	-- STA @3                  	; armazena 0 no milhar
tmp(72)	:= "0001000000100";	-- LDA @4                  	; carrega o valor atual da dezena de milhar
tmp(73)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da dezena de milhar
tmp(74)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(75)	:= "0111001001110";	-- JEQ .INCREMENTA_CMILHAR 	; se for, incrementa a centena de milhar
tmp(76)	:= "0101000000100";	-- STA @4                  	; armazena o novo valor da dezena de milhar
tmp(77)	:= "0110000101101";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(78)	:= "0100000000000";	-- LDI $0                  	; carrega 0
tmp(79)	:= "0101000000100";	-- STA @4                  	; armazena 0 na dezena de milhar
tmp(80)	:= "0001000000101";	-- LDA @5                  	; carrega o valor atual da centena de milhar
tmp(81)	:= "0010000000110";	-- ADD @6                  	; incrementa o valor da centena de milhar
tmp(82)	:= "1000000000111";	-- CEQ @7                  	; verifica se é igual a 10
tmp(83)	:= "0111001010110";	-- JEQ .INCREMENTA_MILHAO  	; se for, zera tudo
tmp(84)	:= "0101000000101";	-- STA @5                  	; armazena o novo valor da centena de milhar
tmp(85)	:= "0110000101101";	-- JMP .FIM_INCREMENTA     	; sai da função
tmp(86)	:= "0100000000000";	-- LDI $0  	; carrega 0
tmp(87)	:= "0101000000101";	-- STA $5  	; armazena 0 na centena de milhar
tmp(88)	:= "0110000101101";	-- JMP .FIM_INCREMENTA
tmp(89)	:= "0001000000000";	-- LDA @0      	; carrega o valor da unidade
tmp(90)	:= "0101100100000";	-- STA @288    	; armazena o 0 no HEX 0
tmp(91)	:= "0001000000001";	-- LDA @1      	; carrega o valor da dezena
tmp(92)	:= "0101100100001";	-- STA @289    	; armazena o 0 no HEX 1
tmp(93)	:= "0001000000010";	-- LDA @2      	; carrega o valor da centena
tmp(94)	:= "0101100100010";	-- STA @290    	; armazena o 0 no HEX 2
tmp(95)	:= "0001000000011";	-- LDA @3      	; carrega o valor do milhar
tmp(96)	:= "0101100100011";	-- STA @291    	; armazena o 0 no HEX 3
tmp(97)	:= "0001000000100";	-- LDA @4      	; carrega o valor da dezena de milhar
tmp(98)	:= "0101100100100";	-- STA @292    	; armazena o 0 no HEX 4
tmp(99)	:= "0001000000101";	-- LDA @5      	; carrega o valor da centena de milhar
tmp(100)	:= "0101100100101";	-- STA @293    	; armazena o 0 no HEX 5
tmp(101)	:= "1000000000000";	-- RET
