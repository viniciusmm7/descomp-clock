tmp(0)	:= "0101111111111";	-- STA @511
tmp(1)	:= "0100000000001";	-- LDI $1
tmp(2)	:= "0101000000001";	-- STA @1
tmp(3)	:= "0000000000000";	-- NOP
tmp(4)	:= "0001101100000";	-- LDA @352
tmp(5)	:= "0101100100000";	-- STA @288
tmp(6)	:= "1011000000001";	-- AND @1
tmp(7)	:= "0101100100001";	-- STA @289
tmp(8)	:= "0000000000000";	-- NOP
tmp(9)	:= "0110000000011";	-- JMP @3
